module cnt(
  input clk,
  input rst_n,
  output clk_1k, 
);


endmodule
