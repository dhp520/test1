module


endmodule
